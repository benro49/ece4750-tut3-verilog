module top;
	initial begin
		$display("Hello world and more!!!");
	end
endmodule
